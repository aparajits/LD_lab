module nand_not(c,a);
input a;
output c;
nand n1(c,a,a);
endmodule
